magic
tech scmos
timestamp 1638804071
<< nwell >>
rect -39 -8 37 26
<< ntransistor >>
rect -21 -51 -18 -42
rect -6 -51 -3 -42
rect 12 -51 15 -42
<< ptransistor >>
rect -21 0 -18 14
rect -6 0 -3 14
rect 12 0 15 14
<< ndiffusion >>
rect -41 -50 -39 -42
rect -31 -50 -21 -42
rect -41 -51 -21 -50
rect -18 -51 -6 -42
rect -3 -51 12 -42
rect 15 -50 19 -42
rect 27 -50 42 -42
rect 15 -51 42 -50
<< pdiffusion >>
rect -23 6 -21 14
rect -31 0 -21 6
rect -18 10 -6 14
rect -18 2 -16 10
rect -8 2 -6 10
rect -18 0 -6 2
rect -3 6 -1 14
rect 7 6 12 14
rect -3 0 12 6
rect 15 6 19 14
rect 15 0 27 6
<< ndcontact >>
rect -39 -50 -31 -42
rect 19 -50 27 -42
<< pdcontact >>
rect -31 6 -23 14
rect -16 2 -8 10
rect -1 6 7 14
rect 19 6 27 14
<< polysilicon >>
rect -21 14 -18 26
rect -6 14 -3 26
rect 12 14 15 26
rect -21 -42 -18 0
rect -6 -42 -3 0
rect 12 -42 15 0
rect -21 -54 -18 -51
rect -6 -54 -3 -51
rect 12 -54 15 -51
<< metal1 >>
rect -46 20 41 24
rect -31 14 -23 20
rect -1 14 8 20
rect -31 5 -23 6
rect -8 2 -7 10
rect 7 6 8 14
rect -16 -12 -7 2
rect 19 -12 27 6
rect -16 -16 77 -12
rect 19 -42 27 -16
rect -39 -57 -31 -50
rect -42 -61 45 -57
<< labels >>
rlabel metal1 -28 22 -28 22 5 vdd
rlabel metal1 -14 -59 -14 -59 1 gnd
<< end >>
