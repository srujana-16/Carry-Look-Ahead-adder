magic
tech scmos
timestamp 1637345551
<< nwell >>
rect -44 12 16 34
rect 37 6 100 37
<< polysilicon >>
rect -27 28 -23 31
rect -6 28 -2 31
rect 59 28 63 34
rect -27 -10 -23 18
rect -24 -15 -23 -10
rect -6 -12 -2 18
rect 59 -10 63 18
rect -27 -26 -23 -15
rect -4 -17 -2 -12
rect -6 -26 -2 -17
rect -27 -40 -23 -34
rect -6 -39 -2 -34
rect 59 -36 63 -17
rect 59 -49 63 -45
<< ndiffusion >>
rect -34 -34 -27 -26
rect -23 -34 -6 -26
rect -2 -34 -1 -26
rect 35 -44 46 -36
rect 54 -44 59 -36
rect 35 -45 59 -44
rect 63 -44 82 -36
rect 90 -44 98 -36
rect 63 -45 98 -44
<< pdiffusion >>
rect -30 20 -27 28
rect -38 18 -27 20
rect -23 20 -18 28
rect -10 20 -6 28
rect -23 18 -6 20
rect -2 20 1 28
rect 9 20 10 28
rect -2 18 10 20
rect 54 20 59 28
rect 46 18 59 20
rect 63 20 82 28
rect 63 18 90 20
<< metal1 >>
rect -38 41 95 49
rect -38 28 -30 41
rect 1 28 9 41
rect 46 28 54 41
rect -18 1 -10 20
rect -18 -6 7 1
rect 3 -10 7 -6
rect -38 -15 -29 -10
rect -24 -15 -22 -10
rect -18 -17 -9 -12
rect -4 -17 -2 -12
rect 3 -17 51 -10
rect 3 -26 7 -17
rect -42 -46 -34 -34
rect 82 -36 90 20
rect -42 -54 14 -46
rect 5 -59 14 -54
rect 46 -59 54 -44
rect 82 -59 90 -44
rect 5 -67 108 -59
<< ntransistor >>
rect -27 -34 -23 -26
rect -6 -34 -2 -26
rect 59 -45 63 -36
<< ptransistor >>
rect -27 18 -23 28
rect -6 18 -2 28
rect 59 18 63 28
<< polycontact >>
rect -29 -15 -24 -10
rect -9 -17 -4 -12
rect 51 -17 63 -10
<< ndcontact >>
rect -42 -34 -34 -26
rect -1 -34 7 -26
rect 46 -44 54 -36
rect 82 -44 90 -36
<< pdcontact >>
rect -38 20 -30 28
rect -18 20 -10 28
rect 1 20 9 28
rect 46 20 54 28
rect 82 20 90 28
<< labels >>
rlabel metal1 -38 -15 -22 -10 1 p
rlabel metal1 -18 -17 -2 -12 1 q
rlabel metal1 23 45 23 45 5 vdd
rlabel metal1 24 -63 24 -63 1 gnd
rlabel metal1 87 -10 87 -10 1 y
<< end >>
