* SPICE3 file created from or4.ext - technology: scmos

.option scale=0.09u

M1000 not_cla_0/a_3_n37# not_cla_0/a_0_n40# not_cla_0/vdd not_cla_0/w_n20_n1# pfet w=9 l=3
+  ad=135 pd=48 as=117 ps=44
M1001 not_cla_0/a_3_n37# not_cla_0/a_0_n40# not_cla_0/gnd Gnd nfet w=9 l=3
+  ad=225 pd=68 as=198 ps=62
M1002 a_n5_9# a_n8_n59# a_n21_9# w_n42_0# pfet w=12 l=3
+  ad=156 pd=50 as=156 ps=50
M1003 gnd a_23_n59# a_11_n56# Gnd nfet w=8 l=3
+  ad=352 pd=136 as=96 ps=40
M1004 a_11_9# a_8_n60# a_n5_9# w_n42_0# pfet w=12 l=3
+  ad=144 pd=48 as=0 ps=0
M1005 gnd a_n8_n59# a_n21_n56# Gnd nfet w=8 l=3
+  ad=0 pd=0 as=104 ps=42
M1006 a_n21_n56# a_n24_n59# gnd Gnd nfet w=8 l=3
+  ad=0 pd=0 as=0 ps=0
M1007 a_n21_9# a_n24_n59# vdd w_n42_0# pfet w=12 l=3
+  ad=0 pd=0 as=120 ps=44
M1008 gnd a_23_n59# a_11_9# w_n42_0# pfet w=12 l=3
+  ad=120 pd=44 as=0 ps=0
M1009 a_11_n56# a_8_n60# gnd Gnd nfet w=8 l=3
+  ad=0 pd=0 as=0 ps=0
C0 not_cla_0/a_3_n37# not_cla_0/gnd 0.09fF
C1 gnd a_n21_n56# 0.05fF
C2 w_n42_0# gnd 0.06fF
C3 gnd a_11_n56# 0.12fF
C4 w_n42_0# a_n24_n59# 0.13fF
C5 not_cla_0/w_n20_n1# not_cla_0/a_0_n40# 0.09fF
C6 w_n42_0# a_n8_n59# 0.13fF
C7 not_cla_0/w_n20_n1# not_cla_0/vdd 0.08fF
C8 w_n42_0# a_8_n60# 0.13fF
C9 not_cla_0/w_n20_n1# not_cla_0/a_3_n37# 0.05fF
C10 not_cla_0/a_0_n40# not_cla_0/vdd 0.08fF
C11 w_n42_0# a_23_n59# 0.13fF
C12 w_n42_0# vdd 0.05fF
C13 not_cla_0/vdd not_cla_0/a_3_n37# 0.06fF
C14 a_11_n56# Gnd 0.02fF
C15 a_n21_n56# Gnd 0.02fF
C16 gnd Gnd 0.79fF
C17 vdd Gnd 0.41fF
C18 a_23_n59# Gnd 0.38fF
C19 a_8_n60# Gnd 0.40fF
C20 a_n8_n59# Gnd 0.39fF
C21 a_n24_n59# Gnd 0.38fF
C22 w_n42_0# Gnd 2.45fF
C23 not_cla_0/gnd Gnd 0.20fF
C24 not_cla_0/a_3_n37# Gnd 0.14fF
C25 not_cla_0/vdd Gnd 0.12fF
C26 not_cla_0/a_0_n40# Gnd 0.26fF
C27 not_cla_0/w_n20_n1# Gnd 0.93fF
