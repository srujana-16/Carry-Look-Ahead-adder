magic
tech scmos
timestamp 1638846014
<< polysilicon >>
rect -138 414 902 429
rect 920 414 937 429
rect -138 396 249 409
rect 259 396 937 409
rect -138 394 937 396
rect -136 385 939 387
rect -136 372 586 385
rect 600 372 939 385
rect -139 364 936 365
rect -139 350 273 364
rect 283 362 936 364
rect 283 350 380 362
rect 387 350 936 362
rect -137 342 938 343
rect -137 328 494 342
rect 511 328 938 342
rect -136 320 939 321
rect -136 306 302 320
rect 312 318 939 320
rect 312 306 395 318
rect 402 306 939 318
rect 414 296 421 297
rect -137 295 938 296
rect -137 293 335 295
rect -137 281 -88 293
rect -72 290 335 293
rect -72 282 152 290
rect 159 282 335 290
rect -72 281 335 282
rect 345 293 938 295
rect 345 281 414 293
rect 421 281 938 293
rect -137 272 938 275
rect -137 260 -112 272
rect -95 260 938 272
rect 382 135 385 137
rect 397 135 400 137
rect 415 135 418 137
rect 593 42 596 67
rect 607 43 610 63
rect 622 42 625 65
rect 247 -12 251 10
rect 274 -14 278 9
rect 304 -14 308 10
rect 336 -13 340 11
rect 874 -103 903 -99
rect 228 -174 231 -159
rect 242 -174 245 -158
rect 257 -174 260 -157
<< polycontact >>
rect 902 414 920 429
rect 249 396 259 410
rect 586 372 600 385
rect 273 350 283 364
rect 380 350 387 362
rect 494 327 511 342
rect 302 306 312 320
rect 395 306 402 318
rect -88 280 -72 293
rect 152 282 159 290
rect 335 281 345 295
rect 414 281 421 293
rect -112 259 -95 272
rect 382 137 386 143
rect 397 137 401 143
rect 415 137 419 143
rect 507 77 511 81
rect 591 67 596 72
rect 605 63 612 70
rect 622 65 627 70
rect 246 10 254 23
rect 271 9 284 28
rect 302 10 315 29
rect 333 11 343 25
rect 681 -2 688 9
rect 903 -105 913 -93
rect 418 -113 426 -105
rect 220 -159 231 -152
rect 235 -158 246 -146
rect 256 -157 267 -145
rect 936 -161 946 -149
rect 312 -209 322 -202
<< metal1 >>
rect 907 392 915 414
rect 383 362 386 363
rect -110 88 -96 259
rect 130 94 138 110
rect 89 92 138 94
rect 89 91 133 92
rect -110 82 -23 88
rect -110 78 -96 82
rect 274 33 283 350
rect 380 346 387 350
rect 273 28 283 33
rect 303 29 312 306
rect 335 182 344 281
rect 382 252 386 346
rect 494 342 509 344
rect 906 332 915 392
rect 395 318 402 320
rect 382 186 385 252
rect 334 177 344 182
rect 194 15 246 17
rect 192 10 246 15
rect 254 10 271 17
rect 192 7 200 10
rect 334 25 343 177
rect 382 143 385 179
rect 397 143 400 306
rect 414 293 421 297
rect 415 143 418 281
rect 494 182 509 327
rect 906 315 914 332
rect 905 298 914 315
rect 493 178 560 182
rect 565 178 588 182
rect 493 176 588 178
rect 683 176 740 181
rect 477 81 483 97
rect 477 77 507 81
rect 522 67 591 72
rect 726 70 733 176
rect 905 149 913 298
rect 905 134 914 149
rect 627 65 733 70
rect 906 67 914 134
rect 905 55 914 67
rect 191 -148 200 7
rect 631 -1 681 9
rect 905 -11 913 55
rect 904 -27 913 -11
rect 369 -104 372 -49
rect 904 -93 912 -27
rect 434 -97 577 -96
rect 434 -98 679 -97
rect 434 -104 689 -98
rect 369 -105 426 -104
rect 472 -105 689 -104
rect 369 -113 418 -105
rect 574 -106 689 -105
rect 369 -114 372 -113
rect 669 -137 689 -106
rect 191 -152 235 -148
rect 191 -158 220 -152
rect 231 -158 235 -152
rect 669 -146 831 -137
rect 669 -147 689 -146
rect 909 -148 919 -147
rect 884 -149 940 -148
rect 687 -160 847 -151
rect 884 -159 936 -149
rect 884 -160 910 -159
rect 915 -160 936 -159
rect 265 -202 276 -200
rect 687 -202 707 -160
rect 935 -161 936 -160
rect 958 -161 993 -149
rect 265 -207 312 -202
rect 274 -209 312 -207
rect 507 -203 707 -202
rect 411 -204 707 -203
rect 333 -211 707 -204
rect 756 -176 861 -167
rect 334 -212 516 -211
rect 756 -212 776 -176
rect 334 -213 439 -212
rect 755 -215 776 -212
rect 755 -312 775 -215
rect 755 -327 776 -312
rect 756 -358 776 -327
rect 378 -366 776 -358
rect 379 -367 776 -366
<< m2contact >>
rect 154 106 159 112
rect -11 79 -6 86
rect 381 179 386 186
rect 560 178 565 185
rect 250 -366 258 -358
rect 272 -368 280 -360
<< metal2 >>
rect -87 86 -75 294
rect 154 112 158 291
rect 250 279 256 410
rect 250 271 257 279
rect 251 188 257 271
rect 588 252 595 385
rect 588 251 750 252
rect 588 245 751 251
rect 250 180 257 188
rect 744 217 751 245
rect 250 156 256 180
rect 386 179 560 185
rect 383 178 560 179
rect 565 178 566 185
rect 290 156 296 157
rect 247 151 296 156
rect -87 79 -11 86
rect -87 78 -6 79
rect -87 77 -75 78
rect 246 45 252 46
rect 290 45 296 151
rect 744 116 752 217
rect 604 109 766 116
rect 605 63 612 109
rect 246 40 296 45
rect 163 20 193 21
rect 246 20 252 40
rect 290 38 296 40
rect 163 14 254 20
rect 163 11 169 14
rect 184 13 254 14
rect 162 -32 169 11
rect 246 9 252 13
rect 162 -152 170 -32
rect 745 -80 752 109
rect 162 -159 232 -152
rect 163 -208 170 -159
rect 744 -207 752 -80
rect 163 -281 171 -208
rect 164 -357 171 -281
rect 423 -237 429 -236
rect 745 -237 752 -207
rect 423 -242 757 -237
rect 423 -297 429 -242
rect 422 -308 429 -297
rect 164 -358 257 -357
rect 164 -365 250 -358
rect 164 -367 171 -365
rect 272 -427 278 -368
rect 271 -428 363 -427
rect 422 -428 428 -308
rect 271 -435 428 -428
rect 354 -436 428 -435
<< metal3 >>
rect 302 15 516 19
rect 303 10 516 15
rect 317 9 516 10
rect 256 -148 405 -147
rect 493 -148 515 9
rect 256 -157 515 -148
rect 399 -158 515 -157
rect 493 -159 515 -158
use and_cla  and_cla_0
timestamp 1638789926
transform 1 0 6 0 1 95
box -44 -67 108 49
use or_cla  or_cla_0
timestamp 1638834781
transform 1 0 156 0 1 110
box -31 -85 114 51
use nand  nand_0
timestamp 1638804071
transform 1 0 403 0 1 109
box -46 -61 77 26
use and_cla  and_cla_1
timestamp 1638789926
transform 1 0 598 0 1 191
box -44 -67 108 49
use not_cla  not_cla_0
timestamp 1638804473
transform 1 0 508 0 1 93
box -23 -44 34 26
use and4  and4_0
timestamp 1638814469
transform 1 0 292 0 1 -59
box -67 -83 164 65
use nor3  nor3_0
timestamp 1638807410
transform 1 0 617 0 1 38
box -39 -69 101 14
use nor3  nor3_1
timestamp 1638807410
transform 1 0 252 0 1 -175
box -39 -69 101 14
use or4  or4_0
timestamp 1638814915
transform 1 0 850 0 1 -133
box -42 -77 126 47
use and_cla  and_cla_2
timestamp 1638789926
transform 1 0 290 0 1 -351
box -44 -67 108 49
<< labels >>
rlabel polysilicon -131 265 -131 265 1 p1
rlabel polysilicon -129 287 -129 287 1 g1
rlabel polysilicon -130 311 -130 311 1 p2
rlabel polysilicon -132 336 -132 336 1 g2
rlabel polysilicon -132 357 -132 357 1 p3
rlabel polysilicon -132 380 -132 380 1 g3
rlabel polysilicon -131 401 -131 401 1 p4
rlabel polysilicon -131 420 -131 420 1 g4
rlabel metal1 91 92 91 92 1 p2g1
rlabel space 524 82 524 82 1 p3p2g1
rlabel space 684 182 684 182 1 p3g2
rlabel metal1 483 -100 483 -100 1 p4p3p2g1
rlabel space 263 96 263 96 1 c2
rlabel space 697 4 697 4 1 c3
rlabel metal1 339 -208 339 -208 1 p4p3g2
rlabel metal1 382 -362 382 -362 1 p4g3
rlabel metal1 986 -156 986 -156 1 cout
<< end >>
