magic
tech scmos
timestamp 1637338390
<< nwell >>
rect -99 29 113 57
<< ntransistor >>
rect -71 -15 -68 -4
rect -20 -13 -17 -2
rect 34 -13 37 -2
rect 84 -12 87 -1
<< ptransistor >>
rect -73 36 -70 51
rect -18 36 -15 51
rect 34 36 37 51
rect 84 36 87 51
<< ndiffusion >>
rect -40 -3 -20 -2
rect -95 -5 -71 -4
rect -95 -13 -87 -5
rect -78 -13 -71 -5
rect -95 -15 -71 -13
rect -68 -5 -45 -4
rect -68 -13 -60 -5
rect -51 -13 -45 -5
rect -40 -11 -35 -3
rect -26 -11 -20 -3
rect -40 -13 -20 -11
rect -17 -4 10 -2
rect -17 -12 -9 -4
rect 0 -12 10 -4
rect -17 -13 10 -12
rect 14 -4 34 -2
rect 14 -12 19 -4
rect 28 -12 34 -4
rect 14 -13 34 -12
rect 37 -3 62 -2
rect 37 -11 40 -3
rect 49 -11 62 -3
rect 37 -13 62 -11
rect 65 -3 84 -1
rect 65 -11 68 -3
rect 77 -11 84 -3
rect 65 -12 84 -11
rect 87 -2 115 -1
rect 87 -10 93 -2
rect 102 -10 115 -2
rect 87 -12 115 -10
rect -68 -15 -45 -13
<< pdiffusion >>
rect -90 47 -73 51
rect -90 39 -87 47
rect -78 39 -73 47
rect -90 36 -73 39
rect -70 48 -45 51
rect -70 40 -60 48
rect -51 40 -45 48
rect -70 36 -45 40
rect -42 48 -18 51
rect -42 40 -35 48
rect -26 40 -18 48
rect -42 36 -18 40
rect -15 48 3 51
rect -15 40 -9 48
rect 0 40 3 48
rect -15 36 3 40
rect 9 48 34 51
rect 9 40 16 48
rect 25 40 34 48
rect 9 36 34 40
rect 37 48 54 51
rect 37 40 40 48
rect 49 40 54 48
rect 37 36 54 40
rect 62 48 84 51
rect 62 40 69 48
rect 78 40 84 48
rect 62 36 84 40
rect 87 48 107 51
rect 87 40 93 48
rect 102 40 107 48
rect 87 36 107 40
<< ndcontact >>
rect -87 -13 -78 -5
rect -60 -13 -51 -5
rect -35 -11 -26 -3
rect -9 -12 0 -4
rect 19 -12 28 -4
rect 40 -11 49 -3
rect 68 -11 77 -3
rect 93 -10 102 -2
<< pdcontact >>
rect -87 39 -78 47
rect -60 40 -51 48
rect -35 40 -26 48
rect -9 40 0 48
rect 16 40 25 48
rect 40 40 49 48
rect 69 40 78 48
rect 93 40 102 48
<< polysilicon >>
rect -110 86 87 96
rect -110 -39 -107 86
rect -73 51 -70 59
rect -18 51 -15 86
rect 34 51 37 59
rect 84 51 87 86
rect -73 15 -70 36
rect -18 28 -15 36
rect 34 24 37 36
rect 26 17 37 24
rect 84 19 87 36
rect -73 12 -17 15
rect -71 -4 -68 0
rect -20 -2 -17 12
rect 34 -2 37 17
rect 86 14 87 19
rect 84 -1 87 14
rect 105 9 106 17
rect 114 9 124 17
rect -71 -39 -68 -15
rect -110 -42 -68 -39
rect -20 -63 -17 -13
rect 34 -16 37 -13
rect 84 -16 87 -12
rect 121 -63 124 9
rect -20 -66 124 -63
<< polycontact >>
rect 18 17 26 24
rect 82 14 86 19
rect 106 9 114 17
<< metal1 >>
rect -60 63 0 71
rect -60 48 -51 63
rect -9 48 0 63
rect -87 -5 -78 39
rect -60 -5 -51 40
rect -35 24 -26 40
rect 16 61 78 71
rect 16 48 25 61
rect 69 48 78 61
rect -9 24 0 40
rect -35 17 18 24
rect 26 17 32 24
rect -35 -3 -26 17
rect -9 -4 0 17
rect 40 -3 49 40
rect 74 14 82 19
rect 93 17 102 40
rect 92 9 106 17
rect 114 9 118 17
rect 93 -2 102 9
rect -87 -45 -78 -13
rect 19 -25 28 -12
rect 40 -25 49 -11
rect 68 -25 77 -11
rect 19 -34 77 -25
rect 40 -45 49 -34
rect -87 -54 49 -45
<< labels >>
rlabel metal1 51 -31 51 -30 1 gnd
rlabel metal1 50 66 50 66 1 vdd
rlabel space 74 14 87 19 1 vb
rlabel polycontact 110 13 110 13 1 vbb
rlabel metal1 45 20 45 20 1 vab
rlabel polysilicon 34 21 34 21 1 va
rlabel metal1 -34 68 -34 68 1 vout
<< end >>
